--=================================================================================================
-- Title       : Auxiliary Package
-- Author      : Alberto Caravantes Arranz
-- Date        : 06/04/2025
--=================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package aux_pkg is

    type natural_array is array(0 to 1) of natural;

end package aux_pkg;

package body aux_pkg is

end package body aux_pkg;
